/*
	MODULE:
		Instruction Decode
*/

module InstructionDecoder
(
	input wire	 		Clock,							// 	Input Clock
	input wire 		Reset,							// 	Reset signal
	
);

endmodule
